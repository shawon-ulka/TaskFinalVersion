//TestBench Generation

module tb_frmt4;//TestBench code start

	reg [7:0] a;
	reg [31:0] b;
	wire  c

endmodule//TestBench code end