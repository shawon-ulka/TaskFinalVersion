`timescale 1ns/1ps
module frmt4(a, b, c);

input a; 
input b; 
output c; 
wire [7:0] a;
wire [31:0] b;
reg  c;

endmodule