// Code Generated from Excel
`timescale 1ns/1ps

module frmt4 (
	input	wire	[7:0]	a,
	input	wire	[31:0]	b,
	output	reg		c
);

endmodule